
// functional_partition

// Just instantiate all the submodules (currently just the register and memory state).

// Project foundation includes

`include "hasim_common.bsh"

// mkFunctionalPartition

// Instantiate the submodules

module [HASIM_MODULE] mkFuncp
    //interface:
         ();
    
endmodule
