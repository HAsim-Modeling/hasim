///////////////////////////////////////////////////////////////////////////////
//                                                                           //
// SMIPS_Interfaces.bsv                                                      //
//                                                                           //
// This is the file we hope will be generated by script to hook up all       //
// links and instantiate the top-level module.                               //
//                                                                           //
// Stuff in this file will be similar to a "linking" phase in software.      //
//                                                                           //
// All components of these interfaces should either be:                      //
// A) Get/Puts                                                               //
// B) Client/Servers                                                         //
//    or                                                          	     //
// C) The original interface                                    	     //
///////////////////////////////////////////////////////////////////////////////

import GetPut::*;
import ClientServer::*;
import RegFile::*;


/************* Functional Partition Interface *************/


interface SMIPS_FunctionalPartition;

  //Original interface
  interface Empty orignal;

  //Links For Timing Partition
  
  interface Server#(Tuple2#(SMIPS_Token, SMIPS_Tick), SMIPS_Token) link_tok;
  interface Server#(Tuple3#(SMIPS_Token, SMIPS_Addr, SMIPS_Tick), Tuple2#(SMIPS_Token, SMIPS_Inst)) link_fet;
  interface Server#(Tuple2#(SMIPS_Token, SMIPS_Tick), Tuple2#(SMIPS_Token, SMIPS_DepInfo)) link_dec;
  interface Server#(Tuple2#(SMIPS_Token, SMIPS_Tick), Tuple2#(SMIPS_Token, SMIPS_InstResult)) link_exe;
  interface Server#(Tuple2#(SMIPS_Token, SMIPS_Tick), SMIPS_Token) link_mem;
  interface Server#(Tuple2#(SMIPS_Token, SMIPS_Tick), SMIPS_Token) link_lco;
  interface Server#(Tuple2#(SMIPS_Token, SMIPS_Tick), SMIPS_Token) link_gco;
  
  interface Put#(SMIPS_Token) link_killToken;
  
  //Links For Memory
  
  interface Client#(MemReq#(SMIPS_Token, SMIPS_Addr, SMIPS_Value), MemResp#(SMIPS_Value)) link_to_dmem;
  interface Client#(SMIPS_Addr, SMIPS_Inst) link_to_imem;
  
  interface Get#(SMIPS_Token) link_commit;
  interface Get#(Tuple2#(SMIPS_Token, SMIPS_Token)) link_killRange;
  
endinterface


/************* Timing Partition Interface *************/

                                //The type parameters come from the original interface
interface SMIPS_TimingPartition#(type tick_T, type command_T);

  //TModule
  interface TModule#(tick_T, command_T) original;
  
  // Links for Functional Partition 
  // (Dual of above)
  
  interface Client#(Tuple2#(SMIPS_Token, SMIPS_Tick), SMIPS_Token) link_tok;
  interface Client#(Tuple3#(SMIPS_Token, SMIPS_Addr, SMIPS_Tick), Tuple2#(SMIPS_Token, SMIPS_Inst)) link_fet;
  interface Client#(Tuple2#(SMIPS_Token, SMIPS_Tick), Tuple2#(SMIPS_Token, SMIPS_DepInfo)) link_dec;
  interface Client#(Tuple2#(SMIPS_Token, SMIPS_Tick), Tuple2#(SMIPS_Token, SMIPS_InstResult)) link_exe;
  interface Client#(Tuple2#(SMIPS_Token, SMIPS_Tick), SMIPS_Token) link_mem;
  interface Client#(Tuple2#(SMIPS_Token, SMIPS_Tick), SMIPS_Token) link_lco;
  interface Client#(Tuple2#(SMIPS_Token, SMIPS_Tick), SMIPS_Token) link_gco;
  
  interface Get#(token_T) link_killToken;
  
endinterface



/************* CPU Interface *************/


interface SMIPS_CPU#(type tick_T, type command_T);

  //TModule
  interface TModule#(tick_T, command_T) original;

  // Links To Memory
  // (Handled by Functional Partition)
  
  interface Client#(MemReq#(SMIPS_Token, SMIPS_Addr, SMIPS_Value), MemResp#(SMIPS_Value)) to_dmem;
  interface Client#(SMIPS_Addr, SMIPS_Inst) to_imem;
  
  interface Get#(SMIPS_Token) commit;
  interface Get#(Tuple2#(SMIPS_Token, SMIPS_Token)) killRange; 

endinterface

