package Primitive(primBitToInteger) where

primitive primBitToInteger :: Bit n -> Integer

