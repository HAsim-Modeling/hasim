`include "asim/provides/low_level_platform_interface.bsh"

module mkSystem#(LowLevelPlatformInterface llpi) ();

endmodule

