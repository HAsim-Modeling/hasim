
typedef TOKEN_INDEX TokIndex;

typedef TOKEN_TIMEP_INFO TIMEP_TokInfo;

typedef TOKEN_FUNCP_INFO FUNCP_TokInfo;

typedef TOKEN_TIMEP_EPOCH TIMEP_Epoch;
typedef TOKEN_TIMEP_SCRATCHPAD TIMEP_Scratchpad;

typedef TOKEN_FUNCP_EPOCH FUNCP_Epoch;
typedef TOKEN_FUNCP_SCRATCHPAD FUNCP_Scratchpad;

typedef TOKEN Token;

typedef ASSERTION_SEVERITY AssertionSeverity;

typedef HASIM_MODULE HASim_Module;
