
//HASim library imports
import hasim_base::*;
import hasim_common::*;

//************* Null Controller **************

// module [HASim_Module] mkController#(TModule#(Command, Response) th) ();
module [HASim_Module] mkController();
   
   
   
endmodule

