
import hasim_common::*;

import hasim_traffic_light_function::*;


module [HASIM_MODULE] mkSystem ();

   let tl <- mk_traffic_light();
  
endmodule
