`include "hasim_common.bsh"

//=============== Null Controller ===============
module [HASim_Module] mkController();
endmodule

