
import hasim_common::*;

import hasim_traffic_light_function::*;


module [HASim_Module] mkSystem ();

   let tl <- mk_traffic_light();
  
endmodule
