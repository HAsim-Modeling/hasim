//
// Copyright (C) 2008 Intel Corporation
//
// This program is free software; you can redistribute it and/or
// modify it under the terms of the GNU General Public License
// as published by the Free Software Foundation; either version 2
// of the License, or (at your option) any later version.
//
// This program is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program; if not, write to the Free Software
// Foundation, Inc., 51 Franklin Street, Fifth Floor, Boston, MA  02110-1301, USA.
//

import FIFO::*;
import GetPut::*;
import Connectable::*;

// Project imports

`include "asim/provides/hasim_common.bsh"
`include "asim/provides/soft_connections.bsh"
`include "asim/provides/common_services.bsh"


// ========================================================================
//
//  Interface idioms
//  
// ========================================================================

//
// All functional interface connections have output buffering sufficient
// for avoiding deadlocks in standard multiplexed models.  The standard
// multiplexed controller allows at most one cycle to be active for each
// context.  One slot is thus sufficient for a machine that is single
// issue.
//

module [CONNECTED_MODULE] mkFUNCPInterfaceServer#(String connectionName)
    // Interface:
    (Connection_Server#(t_REQ, t_RSP))
    provisos (Bits#(t_REQ, t_REQ_SZ),
              Bits#(t_RSP, t_RSP_SZ));
     
    CONNECTION_SERVER#(t_REQ, t_RSP) con <- mkConnectionServer(connectionName);

    //
    // Debugging:  track the number of requests to a server that are in
    //             flight.  This is often a good way to debug deadlocks.
    //
    COUNTER#(8) nInFlight <- mkLCounter(0);

    DEBUG_SCAN_FIELD_LIST dbg_list = List::nil;
    dbg_list <- addDebugScanField(dbg_list, "Requests in flight", nInFlight.value);
    let dbgNode <- mkDebugScanNode("FUNCP REGMGR Service: " + connectionName, dbg_list);


    method Bool   reqNotEmpty() = con.reqNotEmpty();
    method t_REQ  getReq() = con.getReq();

    method Action deq();
        con.deq();
        nInFlight.up();
    endmethod


    method Action makeResp(t_RSP data);
        con.makeRsp(data);
        nInFlight.down();
    endmethod

    method Bool   respNotFull() = con.rspNotFull();
endmodule


// ========================================================================
//
//  Global types
//
// ========================================================================

// UP_TO_TWO

typedef union tagged
{
    a ONE;
    Tuple2#(a, a) TWO;
}
    UP_TO_TWO#(parameter type a)
        deriving (Eq, Bits);

function a getFirst(UP_TO_TWO#(a) d);

    case (d) matches
        tagged ONE .x:         return x;
        tagged TWO {.x1, .x2}: return x1;
    endcase

endfunction

function Bool hasSecond(UP_TO_TWO#(a) d);

    case (d) matches
        tagged ONE .x:         return False;
        tagged TWO {.x1, .x2}: return True;
    endcase

endfunction

function Maybe#(a) getSecond(UP_TO_TWO#(a) d);

    case (d) matches
        tagged ONE .x:         return tagged Invalid;
        tagged TWO {.x1, .x2}: return tagged Valid x2;
    endcase

endfunction

function a getSecondOfTwo(UP_TO_TWO#(a) d);

    case (d) matches
        tagged ONE .x:         return ?;
        tagged TWO {.x1, .x2}: return x2;
    endcase

endfunction


//
// Destination registers.  Architectural and physical registers are kept in
// separate lists because some slots get a physical register even when no
// architectural register is allocated.  (E.g. store data.)
//

typedef struct
{
    Vector#(ISA_MAX_DSTS, Maybe#(ISA_REG_INDEX)) ar;
    ISA_INST_DSTS pr;
}
REGMGR_DST_REGS
    deriving (Bits, Eq);
