
//HASim library imports
import HASim::*;

//HASim model-specific imports
import ISA::*;

//************* Null Controller **************

module [HASim_Module] mkController#(TModule#(Command, Response) th) ();
   
   
   
endmodule

