import soft_connections::*;

typedef Connected_Module HASim_Module;
