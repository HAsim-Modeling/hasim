import GetPut::*;
import RegFile::*;
import FIFO::*;
import Vector::*;

import Interfaces::*;
import Primitive::*;
import ValueVector::*;

