
//HASim library imports
import HASim::*;

//HASim model-specific imports
import NullISA::*;

//************* Null Controller **************

module [HASim_Module] mkController#(TModule#(Command, Response) th) ();
   
   
   
endmodule

