
interface TopLevelWires;
endinterface

module mkTopLevelWires (TopLevelWires);
endmodule
