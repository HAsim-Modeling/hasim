import bluespec_common::*;
import bluespec_system::*;

(* synthesize *)
module mkModel();

    let system <- mkSystem();

endmodule

