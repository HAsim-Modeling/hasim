import hasim_common::*;
import dme_alg::*;

module [HASim_Module] mkSystem ();
   
  let alg <- mkDME_Alg();
  
endmodule
