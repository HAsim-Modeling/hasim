import hasim_common::*;
import afu_alg::*;

module [HASim_Module] mkSystem ();
   
  let alg <- mkAFU_Alg();
  
endmodule
