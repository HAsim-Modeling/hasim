import soft_connections::*;

typedef Connected_Module HASIM_MODULE;
