typedef Bit#(1) UNIT;
