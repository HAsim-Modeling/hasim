import FIFO::*;

import hasim_common::*;
import soft_connections::*;

/* -------------------------------------------------------------------------- */
// The StallPorts model a ping-pong buffer/double buffer.
//
// Description of a ping-pong buffer
// A ping-pong buffer is an implementation of a pipeline latch which has
// storage for two cycles worth of information. If at the beginning of a cycle,
// both entries in the buffer are occupied, the producer will not do any work,
// regardless of whether the consumer plans to consume an entry in that cycle.
// The advantage of this implementation is that there is no combinational path
// from the consumer to the producer. For those familiar with bluespec, this is
// exactly the bluespec mkFIFO.
//
// Here is an example that demonstrates the operation of a ping pong buffer as
// well as bubble squishing. A-F are instructions, FDXMW are pipeline stages.
// || is the ping-pong buffer and S represents a stall. Note that unlike
// conventional pipeline diagrams, I am showing the instructions as sitting
// inside the buffer as opposed to inside a stage.
//
// time       F  ||  D  ||  X  ||  M  ||  W
//    0
//    1           A
//    2           B      A
//    3           C      B      A  S            # S = stall due to cache-miss
//    4           D      C     BA  S
//    5           E     DC     BA
//    6          FE     DC      B      A
//    7          FE  S1  D      C      B        # S1 = stall due to dependency on B
//    8          FE  S1         D  S2  C        # S2 = stall due to cache miss
//    9          FE             D  S2
//   10           F      E      D  S2           # bubble squished
//

/* -------------------------------------------------------------------------- */
// StallPorts Interface:
//
// StallPorts guard the producer from enq-ing valid data when the modelled
// buffering is fully occupied. Only when canSend is True, the producer can
// _send_ valid data. When canSend is False, the producer must _pass_ instead.
// A pass is equivalent to a send-Invalid, but can only be called when the
// buffers are full. A producer must perform exactly one of the following
// actions every model cycle: (a) send valid data, (b) send invalid, or (c)
// pass.
//
// The consumer side can choose to either receive data for a cycle, or pass.
// Since a module may wish to base this decision on the contents of the first
// entry in the buffer, there is also a peek method which will show the data
// without removing it from the buffer. The receive method, on the other hand,
// and also deq it from the fifo.

/* -------------------------------------------------------------------------- */
// Implementation Notes:
//
// The pC & cC are state for a 4 stage FSM as shown:
//
// State pC  cC        Description                       Action
//   A    0   0  Beginning of model cycle     None.
//   B    0   1  Consumer model cycle ended   Block consumer from consuming more data.
//   C    1   0  Producer model cycle ended   Block producer from producing more data.
//   D    1   1  Both P&C model cycles ended  Determine canSend & canReceive for next cycle.
//
// Legal paths: A -> B -> D -> A and A -> C -> D -> A
//
// Note that the implementation allows the producer and consumer to "finish"
// their model cycle in any order, but prevents them from going ahead for more
// than 1 model cycle.

interface PORT_STALL_SEND#(type a);
    method Action doEnq(a x);
    method Action noEnq();
    method Bool   canEnq();
    interface INSTANCE_CONTROL_IN_OUT#(1) ctrl;

endinterface

interface PORT_STALL_RECV#(type a);
    method Action noDeq();
    method Action doDeq();
    method ActionValue#(Maybe#(a)) receive();
    interface INSTANCE_CONTROL_IN_OUT#(1) ctrl;
endinterface


interface PORT_STALL_SEND_MULTIPLEXED#(type ni, type a);
    method Action doEnq(INSTANCE_ID#(ni) iid, a x);
    method Action noEnq(INSTANCE_ID#(ni) iid);
    method Bool   canEnq(INSTANCE_ID#(ni) iid);
    interface INSTANCE_CONTROL_IN_OUT#(ni) ctrl;

endinterface

interface PORT_STALL_RECV_MULTIPLEXED#(type ni, type a);
    method Action noDeq(INSTANCE_ID#(ni) iid);
    method Action doDeq(INSTANCE_ID#(ni) iid);
    method ActionValue#(Maybe#(a)) receive(INSTANCE_ID#(ni) iid);
    interface INSTANCE_CONTROL_IN_OUT#(ni) ctrl;
endinterface


module [HASIM_MODULE] mkPortStallSend#(String s)
                       (PORT_STALL_SEND#(a))
            provisos (Bits#(a, sa),
                      Transmittable#(Maybe#(a)));

    Connection_Receive#(Bool) creditFromQueue <- mkConnectionRecvUG(s + "__cred");

    PORT_SEND#(a) enqToQueue <- mkPortSend(s + "__portDataEnq");

    Reg#(Bool) initCredit <- mkReg(True);

    method Action doEnq (a x) if (initCredit || creditFromQueue.notEmpty());
        if (!initCredit)
        begin
            creditFromQueue.deq();
        end
        initCredit <= False;
        enqToQueue.send(tagged Valid x);
    endmethod

    method Action noEnq() if (initCredit || creditFromQueue.notEmpty());
        if (!initCredit)
        begin
            creditFromQueue.deq();
        end
        initCredit <= False;
        enqToQueue.send(tagged Invalid);
    endmethod

    method Bool canEnq() if (initCredit || creditFromQueue.notEmpty()) = initCredit ? True : creditFromQueue.receive();

    interface INSTANCE_CONTROL_IN_OUT ctrl;

        interface INSTANCE_CONTROL_IN in;
        
            method Bool empty() = !(creditFromQueue.notEmpty() || initCredit); // This is that we have a credit token.
            method Bool balanced() = True;
            method Bool light() = False;
            
            method Maybe#(INSTANCE_ID#(1)) nextReadyInstance() = tagged Valid (?);
            method Action drop() if (initCredit || creditFromQueue.notEmpty());

                if (!initCredit)
                begin
                    creditFromQueue.deq();
                end
                initCredit <= False;
                // Note: we purposely don't write enqToQueue here, since it's a drop.
            
            endmethod
        
        endinterface
        
        interface INSTANCE_CONTROL_OUT out;
            
            method Bool full() = enqToQueue.ctrl.full(); // This is if the output port is full.
            method Bool balanced() = True;
            method Bool heavy() = False;
        
        endinterface

    endinterface

endmodule

module [HASIM_MODULE] mkPortStallRecv#(String s)
        (PORT_STALL_RECV#(a))
            provisos (Bits#(a, sa),
                      Transmittable#(Maybe#(a)));

    Connection_Send#(Bool) creditToProducer <- mkConnectionSendUG(s + "__cred");

    PORT_RECV#(a) enqFromProducer <- mkPortRecv_L0(s + "__portDataEnq");

    FIFOF#(a) fifo <- mkUGSizedFIFOF(2);

    Reg#(Bool) producerCompleted <- mkReg(False); // producer model cycle completed
    Reg#(Bool) consumerCompleted <- mkReg(False); // consumer model cycle completed

    rule endModelCycle (producerCompleted && consumerCompleted && creditToProducer.notFull());

        creditToProducer.send(fifo.notFull());
        producerCompleted <= False;
        consumerCompleted <= False;
        
    endrule

    rule processProducer (!producerCompleted && !enqFromProducer.ctrl.empty() && creditToProducer.notFull());

        let m_val <- enqFromProducer.receive();

        if (m_val matches tagged Valid .val)
        begin
            fifo.enq(val);
        end
        producerCompleted <= True;

    endrule
    
    // NOTE: These depend on higher-level guard checking by local controller
    //       and the consumer module.
    //       !ctrl.empty -> canDeq ? 
    //                          (peek* -> (doDeq | noDeq)) :
    //                          noDeq

    method Action doDeq() if (!consumerCompleted);
        fifo.deq();
        consumerCompleted <= True;
    endmethod

    method ActionValue#(Maybe#(a)) receive() if (!consumerCompleted);
        return fifo.notEmpty() ? tagged Valid fifo.first() : tagged Invalid;
    endmethod

    method Action noDeq() if (!consumerCompleted);
        consumerCompleted <= True;
    endmethod

    interface INSTANCE_CONTROL_IN_OUT ctrl;

        interface INSTANCE_CONTROL_IN in;

            method Bool empty() = consumerCompleted; // This is that we calculated the next state of the FIFO.
            method Bool balanced() = True;
            method Bool light() = False;
            
            method Maybe#(INSTANCE_ID#(ni)) nextReadyInstance() = tagged Valid (?);
            method Action drop();
                consumerCompleted <= True;
            endmethod
        
        endinterface
    
        interface INSTANCE_CONTROL_OUT out;
    
            method Bool full() = !creditToProducer.notFull(); // This is that the credit port is full.
            method Bool balanced() = True;
            method Bool heavy() = False;
        
        endinterface

    endinterface

endmodule


module [HASIM_MODULE] mkPortStallSend_Multiplexed#(String s)
                       (PORT_STALL_SEND_MULTIPLEXED#(ni, a))
            provisos (Bits#(a, sa),
                      Transmittable#(Tuple2#(INSTANCE_ID#(ni), Bool)),
                      Transmittable#(Tuple2#(INSTANCE_ID#(ni), Maybe#(a))));

    Connection_Receive#(Tuple2#(INSTANCE_ID#(ni), Bool)) creditFromQueue <- mkConnectionRecvUG(s + "__cred");

    Connection_Send#(Tuple2#(INSTANCE_ID#(ni), Maybe#(a))) enqToQueue <- mkConnection_Send(s + "__portDataEnq");

    Reg#(Maybe#(INSTANCE_ID#(ni))) initCredit <- mkReg(tagged Valid 0);

    method Action doEnq (INSTANCE_ID#(ni) iid, a x) if (isValid(initCredit) || creditFromQueue.notEmpty());

        if (initCredit matches tagged Valid .cur_iid)
        begin
            if (cur_iid == maxBound)
                initCredit <= tagged Invalid;
            else
                initCredit <= tagged Valid (cur_iid + 1);
        end
        else
        begin
            creditFromQueue.deq();
        end
        
        enqToQueue.send(tuple2(iid, tagged Valid x));

    endmethod

    method Action noEnq(INSTANCE_ID#(ni) iid) if (isValid(initCredit) || creditFromQueue.notEmpty());
        if (initCredit matches tagged Valid .cur_iid)
        begin
            if (cur_iid == maxBound)
                initCredit <= tagged Invalid;
            else
                initCredit <= tagged Valid (cur_iid + 1);
        end
        else
        begin
            creditFromQueue.deq();
        end
        
        enqToQueue.send(tuple2(iid, tagged Invalid));

    endmethod

    method Bool canEnq(INSTANCE_ID#(ni) iid) if (isValid(initCredit) || creditFromQueue.notEmpty());

        if (initCredit matches tagged Invalid)
        begin

            match {.*, .b} = creditFromQueue.receive();
            return b;

        end
        else
        begin

            return True;

        end

    endmethod

    interface INSTANCE_CONTROL_IN_OUT ctrl;

        interface INSTANCE_CONTROL_IN in;
        
            method Bool empty() = !(creditFromQueue.notEmpty() || isValid(initCredit)); // This is that we have a credit token.
            method Bool balanced() = True;
            method Bool light() = False;
            
            method Maybe#(INSTANCE_ID#(ni)) nextReadyInstance();
                if (initCredit matches tagged Valid .iid)
                begin
                    return tagged Valid iid;
                end
                else if (creditFromQueue.notEmpty())
                begin
                    match {.iid, .*} = creditFromQueue.receive();
                    return tagged Valid iid;
                end
                else
                begin
                    return tagged Invalid;
                end
            endmethod

            method Action drop() if (isValid(initCredit) || creditFromQueue.notEmpty());

                if (initCredit matches tagged Valid .cur_iid)
                begin
                    if (cur_iid == maxBound)
                        initCredit <= tagged Invalid;
                    else
                        initCredit <= tagged Valid (cur_iid + 1);
                end
                else
                begin
                    creditFromQueue.deq();
                end

                // Note: we purposely don't write enqToQueue here, since it's a drop.
                
            endmethod
        
        endinterface
        
        interface INSTANCE_CONTROL_OUT out;
            
            method Bool full() = !enqToQueue.notFull(); // This is if the output port is full.
            method Bool balanced() = True;
            method Bool heavy() = False;
        
        endinterface

    endinterface


  
endmodule

module [HASIM_MODULE] mkPortStallRecv_Multiplexed#(String s)
        (PORT_STALL_RECV_MULTIPLEXED#(ni, a))
            provisos (Bits#(a, sa),
                      Transmittable#(Tuple2#(INSTANCE_ID#(ni), Bool)),
                      Transmittable#(Tuple2#(INSTANCE_ID#(ni), Maybe#(a))));

    Connection_Send#(Tuple2#(INSTANCE_ID#(ni), Bool)) creditToProducer <- mkConnectionSendUG(s + "__cred");

    Connection_Receive#(Tuple2#(INSTANCE_ID#(ni), Maybe#(a))) enqFromProducer <- mkConnection_Receive(s + "__portDataEnq");

    // We use these like soft connections which are self-contained.
    FIFOF#(Tuple2#(INSTANCE_ID#(ni), Maybe#(a))) firstQ <- mkFIFOF();
    FIFOF#(Bool) deqQ   <- mkFIFOF();
    FIFOF#(INSTANCE_ID#(ni)) writesQ   <- mkFIFOF();

    Vector#(ni, FIFOF#(a)) fifos <- replicateM(mkUGSizedFIFOF(2));

    rule stage1_enqAndFirst (True);

        match {.iid, .m_enq} = enqFromProducer.receive();
        enqFromProducer.deq();
        
        if (m_enq matches tagged Valid .val)
        begin
            fifos[iid].enq(val);
        end

        if (fifos[iid].notEmpty())
        begin
            firstQ.enq(tuple2(iid, tagged Valid fifos[iid].first()));
        end
        else
        begin
            firstQ.enq(tuple2(iid, tagged Invalid));
        end
        
        writesQ.enq(iid);
        
    endrule

    rule stage2_deqAndCredit (creditToProducer.notFull());

        let iid = writesQ.first();
        writesQ.deq();
 
        if (deqQ.first())
        begin
            fifos[iid].deq();
        end
        deqQ.deq();
        
        creditToProducer.send(tuple2(iid, (fifos[iid].notFull || deqQ.first())));

    endrule
    
    // NOTE: These depend on higher-level guard checking by local controller
    //       and the consumer module.
    //       !ctrl.empty -> canDeq ? 
    //                          (peek* -> (doDeq | noDeq)) :
    //                          noDeq

    method Action doDeq(INSTANCE_ID#(ni) iid);
        deqQ.enq(True);
    endmethod

    method ActionValue#(Maybe#(a)) receive(INSTANCE_ID#(ni) iid);
        match {.iid2, .m_val} = firstQ.first();
        firstQ.deq();
        return m_val; 
    endmethod

    method Action noDeq(INSTANCE_ID#(ni) iid);
        deqQ.enq(False);
    endmethod

    interface INSTANCE_CONTROL_IN_OUT ctrl;

        interface INSTANCE_CONTROL_IN in;

            method Bool empty() = !firstQ.notEmpty();
            method Bool balanced() = True;
            method Bool light() = False;
            method Maybe#(INSTANCE_ID#(ni)) nextReadyInstance();
            
                if (firstQ.notEmpty())
                begin
                    match {.iid, .*} = firstQ.first();
                    return tagged Valid iid;
                end
                else
                begin
                    return tagged Invalid;
                end
            
            endmethod
            
            method Action drop();
                firstQ.deq();
            endmethod
        
        endinterface
    
        interface INSTANCE_CONTROL_OUT out;
    
            method Bool full() = !deqQ.notFull();
            method Bool balanced() = True;
            method Bool heavy() = False;
        
        endinterface

    endinterface



endmodule
